/home/kheyse/private/experiments/regExPE/design/top_genericblock.vhd