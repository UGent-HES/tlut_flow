../rom.vhd