/home/kheyse/private/experiments/regExPE/design/test.vhd