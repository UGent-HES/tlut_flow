../../../../exorw32.vhd