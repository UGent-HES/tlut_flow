/home/kheyse/private/experiments/regExPE/design/counter.vhd