/home/kheyse/private/experiments/regExPE/design/countDecoder.vhd