../../../../treeMult4b.vhd